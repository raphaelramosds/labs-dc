library verilog;
use verilog.vl_types.all;
entity and_gate_vlg_vec_tst is
end and_gate_vlg_vec_tst;
