library verilog;
use verilog.vl_types.all;
entity mux4x1_behavioral_description_vlg_check_tst is
    port(
        S               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end mux4x1_behavioral_description_vlg_check_tst;
