entity ones_counter is
	port(
		A, B, C : in bit;
		S1, S2 : out bit;
	);
end entity;

architecture