ENTITY DigitalClock IS
  PORT (
     : IN BIT;
     : OUT BIT
  );
END;

ARCHITECTURE main OF DigitalClock IS

BEGIN

END;