library verilog;
use verilog.vl_types.all;
entity Mux4x1BehavioralDescription_vlg_check_tst is
    port(
        S               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Mux4x1BehavioralDescription_vlg_check_tst;
