library verilog;
use verilog.vl_types.all;
entity properties_vlg_vec_tst is
end properties_vlg_vec_tst;
