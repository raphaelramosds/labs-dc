library verilog;
use verilog.vl_types.all;
entity and_gate_vlg_check_tst is
    port(
        s               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end and_gate_vlg_check_tst;
