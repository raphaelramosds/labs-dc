library verilog;
use verilog.vl_types.all;
entity ones_counter_vlg_vec_tst is
end ones_counter_vlg_vec_tst;
