ENTITY decoder_for_seven_segment_display IS
	PORT(
		A3, A2, A1, A0: IN BIT;
		S6, S5, S4, S3, S2, S1, S0 : OUT BIT
	);
END;

ARCHITECTURE behav OF decoder_for_seven_segment_display IS
	BEGIN
		S0 <= (A3 AND A2) OR (A3 AND A1) OR (A2 AND NOT(A1) AND NOT(A0)) OR (NOT(A3) AND NOT(A2) AND NOT(A0) AND A1);
		S1 <= (A3 AND A2) OR (A3 AND A1) OR (A2 AND NOT(A1) AND A0) OR (A2 AND A1 AND NOT(A0));
		S2 <= (A3 AND A2) OR (A3 AND A1) OR (NOT(A2) AND A1 AND NOT(A0));
		S3 <= (A3 AND A2) OR (A3 AND A1) OR (A2 AND NOT(A1) AND NOT(A0)) OR (A2 AND A1 AND A0) OR (NOT(A3) AND NOT(A2) AND NOT(A1) AND A0);
		S4 <= A0 OR (A2 AND NOT(A0)) OR (A3 AND A1);
		S5 <= (A3 AND A2) OR (A1 AND A0) OR (A3 AND A1) OR (NOT(A2) AND A1) OR (NOT(A3) AND NOT(A2) AND A0);
		S6 <= (A3 AND A2) OR (A3 AND A1) OR (NOT(A3) AND NOT(A2) AND NOT(A1)) OR (A2 AND A1 AND A0);
END;