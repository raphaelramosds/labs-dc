library verilog;
use verilog.vl_types.all;
entity or_gate_vlg_vec_tst is
end or_gate_vlg_vec_tst;
