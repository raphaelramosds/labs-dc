library verilog;
use verilog.vl_types.all;
entity ones_counter_vlg_check_tst is
    port(
        S1              : in     vl_logic;
        S2              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end ones_counter_vlg_check_tst;
